module vlogger

interface Loggable {
	fields() []Field
}
