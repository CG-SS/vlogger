module vlogger

enum PrimitiveType as u8 {
	bool
	string
	i8
	u8
	i16
	u16
	int
	u32
	i64
	u64
	rune
	f32
	f64
	array
	map
	strut
	error
}