module vlogger

enum Level {
	trace
	debug
	info
	warn
	error
	fatal
	panic
}
