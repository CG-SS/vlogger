module vlogger

pub interface Loggable {
	fields() []Field
}
