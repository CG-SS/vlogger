module vlogger

pub enum PrimitiveType as u8 {
	bool
	string
	i8
	u8
	i16
	u16
	i32
	u32
	i64
	u64
	rune
	f32
	f64
	array
	map
	strut
	error
}
