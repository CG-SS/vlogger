module main

enum TimestampType {
	rfc3339
	rfc3339_nano
	ss
	ss_milli
	ss_micro
	ss_nano
	unix_time
	unix_time_micro
	unix_time_milli
	unix_time_nano
}
