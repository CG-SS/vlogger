module vlogger

fn nop_message_writer(_ Message) {}
